<script>
s
</script>